module SGSR(CLK, GSR);
    input CLK;
    input GSR;
endmodule