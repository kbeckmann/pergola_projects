module OB(I, O);
    input I;
    output O;
    assign O = I;
endmodule