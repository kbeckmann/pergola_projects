module IB(I, O);
    input I;
    output O;
    assign O = I;
endmodule