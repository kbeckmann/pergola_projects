module FD1S3AX(CK, D, Q);

parameter GSR;


    input CK;
    input D;
    output Q;
endmodule